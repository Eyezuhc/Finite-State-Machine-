module thunderbird_wrapper(
    input clk,
    input reset,
    input left,
    input right,
    output [5:0] LED
);
    
endmodule